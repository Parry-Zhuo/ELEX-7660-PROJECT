// ELEX 7660
// File: waveGen.sv
// Description: Determines which data to send to DAC based on input parameters.
// Author: Bryce Reid    Student ID: A01298718    Date: 2025-03-18

module waveGen ( input logic reset_n,   			// reset 
		 input logic wclk,				// wave clock
		 input logic s2,   				// S2 push button
		 input logic [2:0] shape,	   		// wave shape selected signal (0-5)
		 input logic [2:0] depth,			// wave depth selected signal (0-4)
		 output logic onOff,				// on/off signal
		 output logic [11:0] data ) ;     		// data to send to DAC

	logic [7:0] index ;			// 8-bit index for data LUT
	logic [0:255][7:0] SnH_index ;		// a LUT with "random" index values for "randomly" selecting a value from sine LUT for the sample & hold function
	logic [7:0] SnH_index_2 ;		// 8-bit index for selecting the next "random" value from the sample & hold index LUT
	logic [11:0] SnH_value ;		// "randomly" selected value from sine LUT for the sample & hold function
	logic [11:0] next_data ;		
	logic [0:255][11:0] dataTable ;		// active data LUT
	logic [0:4][11:0] sqr_high ;		// for implementing square wave
	logic [0:4][11:0] sqr_low ;		// for implementing square wave

	// assign data LUT for waveform output based on selected shape and depth
	always_comb begin
		case ( { shape, depth } )
			// shape: sine // depth: 1 // OR // // shape: sample & hold // depth: 1 //
			{ 3'd0, 3'd0 }, { 3'd5, 3'd0 } : dataTable = { 12'd2048, 12'd2058, 12'd2068, 12'd2078, 12'd2088, 12'd2098, 12'd2108, 12'd2118, 12'd2127, 12'd2137, 12'd2147, 12'd2157, 12'd2166, 12'd2176, 12'd2185, 12'd2195, 12'd2204, 12'd2213, 12'd2223, 12'd2232, 12'd2241, 12'd2249, 12'd2258, 12'd2267, 12'd2275, 12'd2283, 12'd2291, 12'd2299, 12'd2307, 12'd2315, 12'd2323, 12'd2330, 12'd2337, 12'd2344, 12'd2351, 12'd2358, 12'd2364, 12'd2370, 12'd2376, 12'd2382, 12'd2388, 12'd2393, 12'd2399, 12'd2404, 12'd2409, 12'd2413, 12'd2418, 12'd2422, 12'd2426, 12'd2430, 12'd2433, 12'd2436, 12'd2439, 12'd2442, 12'd2445, 12'd2447, 12'd2449, 12'd2451, 12'd2453, 12'd2454, 12'd2455, 12'd2456, 12'd2457, 12'd2457, 12'd2457, 12'd2457, 12'd2457, 12'd2456, 12'd2455, 12'd2454, 12'd2453, 12'd2451, 12'd2449, 12'd2447, 12'd2445, 12'd2442, 12'd2439, 12'd2436, 12'd2433, 12'd2430, 12'd2426, 12'd2422, 12'd2418, 12'd2413, 12'd2409, 12'd2404, 12'd2399, 12'd2393, 12'd2388, 12'd2382, 12'd2376, 12'd2370, 12'd2364, 12'd2358, 12'd2351, 12'd2344, 12'd2337, 12'd2330, 12'd2323, 12'd2315, 12'd2307, 12'd2299, 12'd2291, 12'd2283, 12'd2275, 12'd2267, 12'd2258, 12'd2249, 12'd2241, 12'd2232, 12'd2223, 12'd2213, 12'd2204, 12'd2195, 12'd2185, 12'd2176, 12'd2166, 12'd2157, 12'd2147, 12'd2137, 12'd2127, 12'd2118, 12'd2108, 12'd2098, 12'd2088, 12'd2078, 12'd2068, 12'd2058, 12'd2048, 12'd2037, 12'd2027, 12'd2017, 12'd2007, 12'd1997, 12'd1987, 12'd1977, 12'd1968, 12'd1958, 12'd1948, 12'd1938, 12'd1929, 12'd1919, 12'd1910, 12'd1900, 12'd1891, 12'd1882, 12'd1872, 12'd1863, 12'd1854, 12'd1846, 12'd1837, 12'd1828, 12'd1820, 12'd1812, 12'd1804, 12'd1796, 12'd1788, 12'd1780, 12'd1772, 12'd1765, 12'd1758, 12'd1751, 12'd1744, 12'd1737, 12'd1731, 12'd1725, 12'd1719, 12'd1713, 12'd1707, 12'd1702, 12'd1696, 12'd1691, 12'd1686, 12'd1682, 12'd1677, 12'd1673, 12'd1669, 12'd1665, 12'd1662, 12'd1659, 12'd1656, 12'd1653, 12'd1650, 12'd1648, 12'd1646, 12'd1644, 12'd1642, 12'd1641, 12'd1640, 12'd1639, 12'd1638, 12'd1638, 12'd1638, 12'd1638, 12'd1638, 12'd1639, 12'd1640, 12'd1641, 12'd1642, 12'd1644, 12'd1646, 12'd1648, 12'd1650, 12'd1653, 12'd1656, 12'd1659, 12'd1662, 12'd1665, 12'd1669, 12'd1673, 12'd1677, 12'd1682, 12'd1686, 12'd1691, 12'd1696, 12'd1702, 12'd1707, 12'd1713, 12'd1719, 12'd1725, 12'd1731, 12'd1737, 12'd1744, 12'd1751, 12'd1758, 12'd1765, 12'd1772, 12'd1780, 12'd1788, 12'd1796, 12'd1804, 12'd1812, 12'd1820, 12'd1828, 12'd1837, 12'd1846, 12'd1854, 12'd1863, 12'd1872, 12'd1882, 12'd1891, 12'd1900, 12'd1910, 12'd1919, 12'd1929, 12'd1938, 12'd1948, 12'd1958, 12'd1968, 12'd1977, 12'd1987, 12'd1997, 12'd2007, 12'd2017, 12'd2027, 12'd2037 } ;
			// shape: sine // depth: 2 // OR // // shape: sample & hold // depth: 2 //
			{ 3'd0, 3'd1 }, { 3'd5, 3'd1 } : dataTable = { 12'd2048, 12'd2068, 12'd2088, 12'd2108, 12'd2128, 12'd2148, 12'd2168, 12'd2188, 12'd2207, 12'd2227, 12'd2247, 12'd2266, 12'd2285, 12'd2304, 12'd2323, 12'd2342, 12'd2361, 12'd2379, 12'd2398, 12'd2416, 12'd2434, 12'd2451, 12'd2469, 12'd2486, 12'd2503, 12'd2519, 12'd2535, 12'd2551, 12'd2567, 12'd2582, 12'd2598, 12'd2612, 12'd2627, 12'd2641, 12'd2654, 12'd2668, 12'd2681, 12'd2693, 12'd2705, 12'd2717, 12'd2728, 12'd2739, 12'd2750, 12'd2760, 12'd2770, 12'd2779, 12'd2788, 12'd2796, 12'd2804, 12'd2812, 12'd2819, 12'd2825, 12'd2831, 12'd2837, 12'd2842, 12'd2847, 12'd2851, 12'd2854, 12'd2858, 12'd2860, 12'd2863, 12'd2864, 12'd2866, 12'd2866, 12'd2866, 12'd2866, 12'd2866, 12'd2864, 12'd2863, 12'd2860, 12'd2858, 12'd2854, 12'd2851, 12'd2847, 12'd2842, 12'd2837, 12'd2831, 12'd2825, 12'd2819, 12'd2812, 12'd2804, 12'd2796, 12'd2788, 12'd2779, 12'd2770, 12'd2760, 12'd2750, 12'd2739, 12'd2728, 12'd2717, 12'd2705, 12'd2693, 12'd2681, 12'd2668, 12'd2654, 12'd2641, 12'd2627, 12'd2612, 12'd2598, 12'd2582, 12'd2567, 12'd2551, 12'd2535, 12'd2519, 12'd2503, 12'd2486, 12'd2469, 12'd2451, 12'd2434, 12'd2416, 12'd2398, 12'd2379, 12'd2361, 12'd2342, 12'd2323, 12'd2304, 12'd2285, 12'd2266, 12'd2247, 12'd2227, 12'd2207, 12'd2188, 12'd2168, 12'd2148, 12'd2128, 12'd2108, 12'd2088, 12'd2068, 12'd2048, 12'd2027, 12'd2007, 12'd1987, 12'd1967, 12'd1947, 12'd1927, 12'd1907, 12'd1888, 12'd1868, 12'd1848, 12'd1829, 12'd1810, 12'd1791, 12'd1772, 12'd1753, 12'd1734, 12'd1716, 12'd1697, 12'd1679, 12'd1661, 12'd1644, 12'd1626, 12'd1609, 12'd1592, 12'd1576, 12'd1560, 12'd1544, 12'd1528, 12'd1513, 12'd1497, 12'd1483, 12'd1468, 12'd1454, 12'd1441, 12'd1427, 12'd1414, 12'd1402, 12'd1390, 12'd1378, 12'd1367, 12'd1356, 12'd1345, 12'd1335, 12'd1325, 12'd1316, 12'd1307, 12'd1299, 12'd1291, 12'd1283, 12'd1276, 12'd1270, 12'd1264, 12'd1258, 12'd1253, 12'd1248, 12'd1244, 12'd1241, 12'd1237, 12'd1235, 12'd1232, 12'd1231, 12'd1229, 12'd1229, 12'd1228, 12'd1229, 12'd1229, 12'd1231, 12'd1232, 12'd1235, 12'd1237, 12'd1241, 12'd1244, 12'd1248, 12'd1253, 12'd1258, 12'd1264, 12'd1270, 12'd1276, 12'd1283, 12'd1291, 12'd1299, 12'd1307, 12'd1316, 12'd1325, 12'd1335, 12'd1345, 12'd1356, 12'd1367, 12'd1378, 12'd1390, 12'd1402, 12'd1414, 12'd1427, 12'd1441, 12'd1454, 12'd1468, 12'd1483, 12'd1497, 12'd1513, 12'd1528, 12'd1544, 12'd1560, 12'd1576, 12'd1592, 12'd1609, 12'd1626, 12'd1644, 12'd1661, 12'd1679, 12'd1697, 12'd1716, 12'd1734, 12'd1753, 12'd1772, 12'd1791, 12'd1810, 12'd1829, 12'd1848, 12'd1868, 12'd1888, 12'd1907, 12'd1927, 12'd1947, 12'd1967, 12'd1987, 12'd2007, 12'd2027 } ;
			// shape: sine // depth: 3 // OR // // shape: sample & hold // depth: 3 //
			{ 3'd0, 3'd2 }, { 3'd5, 3'd2 } : dataTable = { 12'd2048, 12'd2078, 12'd2108, 12'd2138, 12'd2168, 12'd2198, 12'd2228, 12'd2258, 12'd2287, 12'd2317, 12'd2346, 12'd2375, 12'd2404, 12'd2433, 12'd2461, 12'd2490, 12'd2518, 12'd2545, 12'd2573, 12'd2600, 12'd2627, 12'd2653, 12'd2679, 12'd2705, 12'd2730, 12'd2755, 12'd2779, 12'd2803, 12'd2827, 12'd2850, 12'd2873, 12'd2895, 12'd2916, 12'd2937, 12'd2958, 12'd2978, 12'd2997, 12'd3016, 12'd3034, 12'd3052, 12'd3069, 12'd3085, 12'd3101, 12'd3116, 12'd3131, 12'd3145, 12'd3158, 12'd3171, 12'd3182, 12'd3194, 12'd3204, 12'd3214, 12'd3223, 12'd3231, 12'd3239, 12'd3246, 12'd3252, 12'd3258, 12'd3263, 12'd3267, 12'd3270, 12'd3273, 12'd3275, 12'd3276, 12'd3276, 12'd3276, 12'd3275, 12'd3273, 12'd3270, 12'd3267, 12'd3263, 12'd3258, 12'd3252, 12'd3246, 12'd3239, 12'd3231, 12'd3223, 12'd3214, 12'd3204, 12'd3194, 12'd3182, 12'd3171, 12'd3158, 12'd3145, 12'd3131, 12'd3116, 12'd3101, 12'd3085, 12'd3069, 12'd3052, 12'd3034, 12'd3016, 12'd2997, 12'd2978, 12'd2958, 12'd2937, 12'd2916, 12'd2895, 12'd2873, 12'd2850, 12'd2827, 12'd2803, 12'd2779, 12'd2755, 12'd2730, 12'd2705, 12'd2679, 12'd2653, 12'd2627, 12'd2600, 12'd2573, 12'd2545, 12'd2518, 12'd2490, 12'd2461, 12'd2433, 12'd2404, 12'd2375, 12'd2346, 12'd2317, 12'd2287, 12'd2258, 12'd2228, 12'd2198, 12'd2168, 12'd2138, 12'd2108, 12'd2078, 12'd2048, 12'd2017, 12'd1987, 12'd1957, 12'd1927, 12'd1897, 12'd1867, 12'd1837, 12'd1808, 12'd1778, 12'd1749, 12'd1720, 12'd1691, 12'd1662, 12'd1634, 12'd1605, 12'd1577, 12'd1550, 12'd1522, 12'd1495, 12'd1468, 12'd1442, 12'd1416, 12'd1390, 12'd1365, 12'd1340, 12'd1316, 12'd1292, 12'd1268, 12'd1245, 12'd1222, 12'd1200, 12'd1179, 12'd1158, 12'd1137, 12'd1117, 12'd1098, 12'd1079, 12'd1061, 12'd1043, 12'd1026, 12'd1010, 12'd994, 12'd979, 12'd964, 12'd950, 12'd937, 12'd924, 12'd913, 12'd901, 12'd891, 12'd881, 12'd872, 12'd864, 12'd856, 12'd849, 12'd843, 12'd837, 12'd832, 12'd828, 12'd825, 12'd822, 12'd820, 12'd819, 12'd819, 12'd819, 12'd820, 12'd822, 12'd825, 12'd828, 12'd832, 12'd837, 12'd843, 12'd849, 12'd856, 12'd864, 12'd872, 12'd881, 12'd891, 12'd901, 12'd913, 12'd924, 12'd937, 12'd950, 12'd964, 12'd979, 12'd994, 12'd1010, 12'd1026, 12'd1043, 12'd1061, 12'd1079, 12'd1098, 12'd1117, 12'd1137, 12'd1158, 12'd1179, 12'd1200, 12'd1222, 12'd1245, 12'd1268, 12'd1292, 12'd1316, 12'd1340, 12'd1365, 12'd1390, 12'd1416, 12'd1442, 12'd1468, 12'd1495, 12'd1522, 12'd1550, 12'd1577, 12'd1605, 12'd1634, 12'd1662, 12'd1691, 12'd1720, 12'd1749, 12'd1778, 12'd1808, 12'd1837, 12'd1867, 12'd1897, 12'd1927, 12'd1957, 12'd1987, 12'd2017 } ;
			// shape: sine // depth: 4 // OR // // shape: sample & hold // depth: 4 //
			{ 3'd0, 3'd3 }, { 3'd5, 3'd3 } : dataTable = { 12'd2048, 12'd2088, 12'd2128, 12'd2168, 12'd2208, 12'd2248, 12'd2288, 12'd2328, 12'd2367, 12'd2406, 12'd2446, 12'd2484, 12'd2523, 12'd2561, 12'd2599, 12'd2637, 12'd2674, 12'd2711, 12'd2748, 12'd2784, 12'd2820, 12'd2855, 12'd2890, 12'd2924, 12'd2958, 12'd2991, 12'd3023, 12'd3055, 12'd3087, 12'd3117, 12'd3148, 12'd3177, 12'd3206, 12'd3234, 12'd3261, 12'd3288, 12'd3314, 12'd3339, 12'd3363, 12'd3387, 12'd3409, 12'd3431, 12'd3452, 12'd3473, 12'd3492, 12'd3511, 12'd3528, 12'd3545, 12'd3561, 12'd3576, 12'd3590, 12'd3603, 12'd3615, 12'd3626, 12'd3636, 12'd3646, 12'd3654, 12'd3661, 12'd3668, 12'd3673, 12'd3678, 12'd3681, 12'd3684, 12'd3685, 12'd3686, 12'd3685, 12'd3684, 12'd3681, 12'd3678, 12'd3673, 12'd3668, 12'd3661, 12'd3654, 12'd3646, 12'd3636, 12'd3626, 12'd3615, 12'd3603, 12'd3590, 12'd3576, 12'd3561, 12'd3545, 12'd3528, 12'd3511, 12'd3492, 12'd3473, 12'd3452, 12'd3431, 12'd3409, 12'd3387, 12'd3363, 12'd3339, 12'd3314, 12'd3288, 12'd3261, 12'd3234, 12'd3206, 12'd3177, 12'd3148, 12'd3117, 12'd3087, 12'd3055, 12'd3023, 12'd2991, 12'd2958, 12'd2924, 12'd2890, 12'd2855, 12'd2820, 12'd2784, 12'd2748, 12'd2711, 12'd2674, 12'd2637, 12'd2599, 12'd2561, 12'd2523, 12'd2484, 12'd2446, 12'd2406, 12'd2367, 12'd2328, 12'd2288, 12'd2248, 12'd2208, 12'd2168, 12'd2128, 12'd2088, 12'd2048, 12'd2007, 12'd1967, 12'd1927, 12'd1887, 12'd1847, 12'd1807, 12'd1767, 12'd1728, 12'd1689, 12'd1649, 12'd1611, 12'd1572, 12'd1534, 12'd1496, 12'd1458, 12'd1421, 12'd1384, 12'd1347, 12'd1311, 12'd1275, 12'd1240, 12'd1205, 12'd1171, 12'd1137, 12'd1104, 12'd1072, 12'd1040, 12'd1008, 12'd978, 12'd947, 12'd918, 12'd889, 12'd861, 12'd834, 12'd807, 12'd781, 12'd756, 12'd732, 12'd708, 12'd686, 12'd664, 12'd643, 12'd622, 12'd603, 12'd584, 12'd567, 12'd550, 12'd534, 12'd519, 12'd505, 12'd492, 12'd480, 12'd469, 12'd459, 12'd449, 12'd441, 12'd434, 12'd427, 12'd422, 12'd417, 12'd414, 12'd411, 12'd410, 12'd410, 12'd410, 12'd411, 12'd414, 12'd417, 12'd422, 12'd427, 12'd434, 12'd441, 12'd449, 12'd459, 12'd469, 12'd480, 12'd492, 12'd505, 12'd519, 12'd534, 12'd550, 12'd567, 12'd584, 12'd603, 12'd622, 12'd643, 12'd664, 12'd686, 12'd708, 12'd732, 12'd756, 12'd781, 12'd807, 12'd834, 12'd861, 12'd889, 12'd918, 12'd947, 12'd978, 12'd1008, 12'd1040, 12'd1072, 12'd1104, 12'd1137, 12'd1171, 12'd1205, 12'd1240, 12'd1275, 12'd1311, 12'd1347, 12'd1384, 12'd1421, 12'd1458, 12'd1496, 12'd1534, 12'd1572, 12'd1611, 12'd1649, 12'd1689, 12'd1728, 12'd1767, 12'd1807, 12'd1847, 12'd1887, 12'd1927, 12'd1967, 12'd2007 } ;
			// shape: sine // depth: 5 // OR // // shape: sample & hold // depth: 5 //
			{ 3'd0, 3'd4 }, { 3'd5, 3'd4 } : dataTable = { 12'd2048, 12'd2098, 12'd2148, 12'd2198, 12'd2248, 12'd2298, 12'd2348, 12'd2398, 12'd2447, 12'd2496, 12'd2545, 12'd2594, 12'd2642, 12'd2690, 12'd2737, 12'd2784, 12'd2831, 12'd2877, 12'd2923, 12'd2968, 12'd3013, 12'd3057, 12'd3100, 12'd3143, 12'd3185, 12'd3226, 12'd3267, 12'd3307, 12'd3346, 12'd3385, 12'd3423, 12'd3459, 12'd3495, 12'd3530, 12'd3565, 12'd3598, 12'd3630, 12'd3662, 12'd3692, 12'd3722, 12'd3750, 12'd3777, 12'd3804, 12'd3829, 12'd3853, 12'd3876, 12'd3898, 12'd3919, 12'd3939, 12'd3958, 12'd3975, 12'd3992, 12'd4007, 12'd4021, 12'd4034, 12'd4045, 12'd4056, 12'd4065, 12'd4073, 12'd4080, 12'd4085, 12'd4089, 12'd4093, 12'd4094, 12'd4095, 12'd4094, 12'd4093, 12'd4089, 12'd4085, 12'd4080, 12'd4073, 12'd4065, 12'd4056, 12'd4045, 12'd4034, 12'd4021, 12'd4007, 12'd3992, 12'd3975, 12'd3958, 12'd3939, 12'd3919, 12'd3898, 12'd3876, 12'd3853, 12'd3829, 12'd3804, 12'd3777, 12'd3750, 12'd3722, 12'd3692, 12'd3662, 12'd3630, 12'd3598, 12'd3565, 12'd3530, 12'd3495, 12'd3459, 12'd3423, 12'd3385, 12'd3346, 12'd3307, 12'd3267, 12'd3226, 12'd3185, 12'd3143, 12'd3100, 12'd3057, 12'd3013, 12'd2968, 12'd2923, 12'd2877, 12'd2831, 12'd2784, 12'd2737, 12'd2690, 12'd2642, 12'd2594, 12'd2545, 12'd2496, 12'd2447, 12'd2398, 12'd2348, 12'd2298, 12'd2248, 12'd2198, 12'd2148, 12'd2098, 12'd2048, 12'd1997, 12'd1947, 12'd1897, 12'd1847, 12'd1797, 12'd1747, 12'd1697, 12'd1648, 12'd1599, 12'd1550, 12'd1501, 12'd1453, 12'd1405, 12'd1358, 12'd1311, 12'd1264, 12'd1218, 12'd1172, 12'd1127, 12'd1082, 12'd1038, 12'd995, 12'd952, 12'd910, 12'd869, 12'd828, 12'd788, 12'd749, 12'd710, 12'd672, 12'd636, 12'd600, 12'd565, 12'd530, 12'd497, 12'd465, 12'd433, 12'd403, 12'd373, 12'd345, 12'd318, 12'd291, 12'd266, 12'd242, 12'd219, 12'd197, 12'd176, 12'd156, 12'd137, 12'd120, 12'd103, 12'd88, 12'd74, 12'd61, 12'd50, 12'd39, 12'd30, 12'd22, 12'd15, 12'd10, 12'd6, 12'd2, 12'd1, 12'd0, 12'd1, 12'd2, 12'd6, 12'd10, 12'd15, 12'd22, 12'd30, 12'd39, 12'd50, 12'd61, 12'd74, 12'd88, 12'd103, 12'd120, 12'd137, 12'd156, 12'd176, 12'd197, 12'd219, 12'd242, 12'd266, 12'd291, 12'd318, 12'd345, 12'd373, 12'd403, 12'd433, 12'd465, 12'd497, 12'd530, 12'd565, 12'd600, 12'd636, 12'd672, 12'd710, 12'd749, 12'd788, 12'd828, 12'd869, 12'd910, 12'd952, 12'd995, 12'd1038, 12'd1082, 12'd1127, 12'd1172, 12'd1218, 12'd1264, 12'd1311, 12'd1358, 12'd1405, 12'd1453, 12'd1501, 12'd1550, 12'd1599, 12'd1648, 12'd1697, 12'd1747, 12'd1797, 12'd1847, 12'd1897, 12'd1947, 12'd1997 } ;
			// shape: triangle // depth: 1 //
			{ 3'd2, 3'd0 } : dataTable = { 12'd1638, 12'd1644, 12'd1651, 12'd1657, 12'd1664, 12'd1670, 12'd1677, 12'd1683, 12'd1690, 12'd1696, 12'd1702, 12'd1709, 12'd1715, 12'd1722, 12'd1728, 12'd1735, 12'd1741, 12'd1748, 12'd1754, 12'd1761, 12'd1767, 12'd1773, 12'd1780, 12'd1786, 12'd1793, 12'd1799, 12'd1806, 12'd1812, 12'd1819, 12'd1825, 12'd1831, 12'd1838, 12'd1844, 12'd1851, 12'd1857, 12'd1864, 12'd1870, 12'd1877, 12'd1883, 12'd1890, 12'd1896, 12'd1902, 12'd1909, 12'd1915, 12'd1922, 12'd1928, 12'd1935, 12'd1941, 12'd1948, 12'd1954, 12'd1960, 12'd1967, 12'd1973, 12'd1980, 12'd1986, 12'd1993, 12'd1999, 12'd2006, 12'd2012, 12'd2018, 12'd2025, 12'd2031, 12'd2038, 12'd2044, 12'd2051, 12'd2057, 12'd2064, 12'd2070, 12'd2077, 12'd2083, 12'd2089, 12'd2096, 12'd2102, 12'd2109, 12'd2115, 12'd2122, 12'd2128, 12'd2135, 12'd2141, 12'd2147, 12'd2154, 12'd2160, 12'd2167, 12'd2173, 12'd2180, 12'd2186, 12'd2193, 12'd2199, 12'd2205, 12'd2212, 12'd2218, 12'd2225, 12'd2231, 12'd2238, 12'd2244, 12'd2251, 12'd2257, 12'd2264, 12'd2270, 12'd2276, 12'd2283, 12'd2289, 12'd2296, 12'd2302, 12'd2309, 12'd2315, 12'd2322, 12'd2328, 12'd2334, 12'd2341, 12'd2347, 12'd2354, 12'd2360, 12'd2367, 12'd2373, 12'd2380, 12'd2386, 12'd2393, 12'd2399, 12'd2405, 12'd2412, 12'd2418, 12'd2425, 12'd2431, 12'd2438, 12'd2444, 12'd2451, 12'd2457, 12'd2457, 12'd2451, 12'd2444, 12'd2438, 12'd2431, 12'd2425, 12'd2418, 12'd2412, 12'd2405, 12'd2399, 12'd2393, 12'd2386, 12'd2380, 12'd2373, 12'd2367, 12'd2360, 12'd2354, 12'd2347, 12'd2341, 12'd2334, 12'd2328, 12'd2322, 12'd2315, 12'd2309, 12'd2302, 12'd2296, 12'd2289, 12'd2283, 12'd2276, 12'd2270, 12'd2264, 12'd2257, 12'd2251, 12'd2244, 12'd2238, 12'd2231, 12'd2225, 12'd2218, 12'd2212, 12'd2205, 12'd2199, 12'd2193, 12'd2186, 12'd2180, 12'd2173, 12'd2167, 12'd2160, 12'd2154, 12'd2147, 12'd2141, 12'd2135, 12'd2128, 12'd2122, 12'd2115, 12'd2109, 12'd2102, 12'd2096, 12'd2089, 12'd2083, 12'd2077, 12'd2070, 12'd2064, 12'd2057, 12'd2051, 12'd2044, 12'd2038, 12'd2031, 12'd2025, 12'd2018, 12'd2012, 12'd2006, 12'd1999, 12'd1993, 12'd1986, 12'd1980, 12'd1973, 12'd1967, 12'd1960, 12'd1954, 12'd1948, 12'd1941, 12'd1935, 12'd1928, 12'd1922, 12'd1915, 12'd1909, 12'd1902, 12'd1896, 12'd1890, 12'd1883, 12'd1877, 12'd1870, 12'd1864, 12'd1857, 12'd1851, 12'd1844, 12'd1838, 12'd1831, 12'd1825, 12'd1819, 12'd1812, 12'd1806, 12'd1799, 12'd1793, 12'd1786, 12'd1780, 12'd1773, 12'd1767, 12'd1761, 12'd1754, 12'd1748, 12'd1741, 12'd1735, 12'd1728, 12'd1722, 12'd1715, 12'd1709, 12'd1702, 12'd1696, 12'd1690, 12'd1683, 12'd1677, 12'd1670, 12'd1664, 12'd1657, 12'd1651, 12'd1644, 12'd1638 } ;
			// shape: triangle // depth: 2 //
			{ 3'd2, 3'd1 } : dataTable = { 12'd1228, 12'd1241, 12'd1254, 12'd1267, 12'd1280, 12'd1293, 12'd1306, 12'd1319, 12'd1332, 12'd1345, 12'd1357, 12'd1370, 12'd1383, 12'd1396, 12'd1409, 12'd1422, 12'd1435, 12'd1448, 12'd1461, 12'd1474, 12'd1486, 12'd1499, 12'd1512, 12'd1525, 12'd1538, 12'd1551, 12'd1564, 12'd1577, 12'd1590, 12'd1603, 12'd1615, 12'd1628, 12'd1641, 12'd1654, 12'd1667, 12'd1680, 12'd1693, 12'd1706, 12'd1719, 12'd1732, 12'd1744, 12'd1757, 12'd1770, 12'd1783, 12'd1796, 12'd1809, 12'd1822, 12'd1835, 12'd1848, 12'd1860, 12'd1873, 12'd1886, 12'd1899, 12'd1912, 12'd1925, 12'd1938, 12'd1951, 12'd1964, 12'd1977, 12'd1989, 12'd2002, 12'd2015, 12'd2028, 12'd2041, 12'd2054, 12'd2067, 12'd2080, 12'd2093, 12'd2106, 12'd2118, 12'd2131, 12'd2144, 12'd2157, 12'd2170, 12'd2183, 12'd2196, 12'd2209, 12'd2222, 12'd2235, 12'd2247, 12'd2260, 12'd2273, 12'd2286, 12'd2299, 12'd2312, 12'd2325, 12'd2338, 12'd2351, 12'd2363, 12'd2376, 12'd2389, 12'd2402, 12'd2415, 12'd2428, 12'd2441, 12'd2454, 12'd2467, 12'd2480, 12'd2492, 12'd2505, 12'd2518, 12'd2531, 12'd2544, 12'd2557, 12'd2570, 12'd2583, 12'd2596, 12'd2609, 12'd2621, 12'd2634, 12'd2647, 12'd2660, 12'd2673, 12'd2686, 12'd2699, 12'd2712, 12'd2725, 12'd2738, 12'd2750, 12'd2763, 12'd2776, 12'd2789, 12'd2802, 12'd2815, 12'd2828, 12'd2841, 12'd2854, 12'd2866, 12'd2866, 12'd2854, 12'd2841, 12'd2828, 12'd2815, 12'd2802, 12'd2789, 12'd2776, 12'd2763, 12'd2750, 12'd2738, 12'd2725, 12'd2712, 12'd2699, 12'd2686, 12'd2673, 12'd2660, 12'd2647, 12'd2634, 12'd2621, 12'd2609, 12'd2596, 12'd2583, 12'd2570, 12'd2557, 12'd2544, 12'd2531, 12'd2518, 12'd2505, 12'd2492, 12'd2480, 12'd2467, 12'd2454, 12'd2441, 12'd2428, 12'd2415, 12'd2402, 12'd2389, 12'd2376, 12'd2363, 12'd2351, 12'd2338, 12'd2325, 12'd2312, 12'd2299, 12'd2286, 12'd2273, 12'd2260, 12'd2247, 12'd2235, 12'd2222, 12'd2209, 12'd2196, 12'd2183, 12'd2170, 12'd2157, 12'd2144, 12'd2131, 12'd2118, 12'd2106, 12'd2093, 12'd2080, 12'd2067, 12'd2054, 12'd2041, 12'd2028, 12'd2015, 12'd2002, 12'd1989, 12'd1977, 12'd1964, 12'd1951, 12'd1938, 12'd1925, 12'd1912, 12'd1899, 12'd1886, 12'd1873, 12'd1860, 12'd1848, 12'd1835, 12'd1822, 12'd1809, 12'd1796, 12'd1783, 12'd1770, 12'd1757, 12'd1744, 12'd1732, 12'd1719, 12'd1706, 12'd1693, 12'd1680, 12'd1667, 12'd1654, 12'd1641, 12'd1628, 12'd1615, 12'd1603, 12'd1590, 12'd1577, 12'd1564, 12'd1551, 12'd1538, 12'd1525, 12'd1512, 12'd1499, 12'd1486, 12'd1474, 12'd1461, 12'd1448, 12'd1435, 12'd1422, 12'd1409, 12'd1396, 12'd1383, 12'd1370, 12'd1357, 12'd1345, 12'd1332, 12'd1319, 12'd1306, 12'd1293, 12'd1280, 12'd1267, 12'd1254, 12'd1241, 12'd1228 } ;
			// shape: triangle // depth: 3 //
			{ 3'd2, 3'd2 } : dataTable = { 12'd819, 12'd838, 12'd858, 12'd877, 12'd896, 12'd916, 12'd935, 12'd954, 12'd974, 12'd993, 12'd1012, 12'd1032, 12'd1051, 12'd1071, 12'd1090, 12'd1109, 12'd1129, 12'd1148, 12'd1167, 12'd1187, 12'd1206, 12'd1225, 12'd1245, 12'd1264, 12'd1283, 12'd1303, 12'd1322, 12'd1341, 12'd1361, 12'd1380, 12'd1399, 12'd1419, 12'd1438, 12'd1457, 12'd1477, 12'd1496, 12'd1515, 12'd1535, 12'd1554, 12'd1574, 12'd1593, 12'd1612, 12'd1632, 12'd1651, 12'd1670, 12'd1690, 12'd1709, 12'd1728, 12'd1748, 12'd1767, 12'd1786, 12'd1806, 12'd1825, 12'd1844, 12'd1864, 12'd1883, 12'd1902, 12'd1922, 12'd1941, 12'd1960, 12'd1980, 12'd1999, 12'd2018, 12'd2038, 12'd2057, 12'd2077, 12'd2096, 12'd2115, 12'd2135, 12'd2154, 12'd2173, 12'd2193, 12'd2212, 12'd2231, 12'd2251, 12'd2270, 12'd2289, 12'd2309, 12'd2328, 12'd2347, 12'd2367, 12'd2386, 12'd2405, 12'd2425, 12'd2444, 12'd2463, 12'd2483, 12'd2502, 12'd2521, 12'd2541, 12'd2560, 12'd2580, 12'd2599, 12'd2618, 12'd2638, 12'd2657, 12'd2676, 12'd2696, 12'd2715, 12'd2734, 12'd2754, 12'd2773, 12'd2792, 12'd2812, 12'd2831, 12'd2850, 12'd2870, 12'd2889, 12'd2908, 12'd2928, 12'd2947, 12'd2966, 12'd2986, 12'd3005, 12'd3024, 12'd3044, 12'd3063, 12'd3083, 12'd3102, 12'd3121, 12'd3141, 12'd3160, 12'd3179, 12'd3199, 12'd3218, 12'd3237, 12'd3257, 12'd3276, 12'd3276, 12'd3257, 12'd3237, 12'd3218, 12'd3199, 12'd3179, 12'd3160, 12'd3141, 12'd3121, 12'd3102, 12'd3083, 12'd3063, 12'd3044, 12'd3024, 12'd3005, 12'd2986, 12'd2966, 12'd2947, 12'd2928, 12'd2908, 12'd2889, 12'd2870, 12'd2850, 12'd2831, 12'd2812, 12'd2792, 12'd2773, 12'd2754, 12'd2734, 12'd2715, 12'd2696, 12'd2676, 12'd2657, 12'd2638, 12'd2618, 12'd2599, 12'd2580, 12'd2560, 12'd2541, 12'd2521, 12'd2502, 12'd2483, 12'd2463, 12'd2444, 12'd2425, 12'd2405, 12'd2386, 12'd2367, 12'd2347, 12'd2328, 12'd2309, 12'd2289, 12'd2270, 12'd2251, 12'd2231, 12'd2212, 12'd2193, 12'd2173, 12'd2154, 12'd2135, 12'd2115, 12'd2096, 12'd2077, 12'd2057, 12'd2038, 12'd2018, 12'd1999, 12'd1980, 12'd1960, 12'd1941, 12'd1922, 12'd1902, 12'd1883, 12'd1864, 12'd1844, 12'd1825, 12'd1806, 12'd1786, 12'd1767, 12'd1748, 12'd1728, 12'd1709, 12'd1690, 12'd1670, 12'd1651, 12'd1632, 12'd1612, 12'd1593, 12'd1574, 12'd1554, 12'd1535, 12'd1515, 12'd1496, 12'd1477, 12'd1457, 12'd1438, 12'd1419, 12'd1399, 12'd1380, 12'd1361, 12'd1341, 12'd1322, 12'd1303, 12'd1283, 12'd1264, 12'd1245, 12'd1225, 12'd1206, 12'd1187, 12'd1167, 12'd1148, 12'd1129, 12'd1109, 12'd1090, 12'd1071, 12'd1051, 12'd1032, 12'd1012, 12'd993, 12'd974, 12'd954, 12'd935, 12'd916, 12'd896, 12'd877, 12'd858, 12'd838, 12'd819 } ;
			// shape: triangle // depth: 4 //
			{ 3'd2, 3'd3 } : dataTable = { 12'd410, 12'd435, 12'd461, 12'd487, 12'd513, 12'd538, 12'd564, 12'd590, 12'd616, 12'd642, 12'd667, 12'd693, 12'd719, 12'd745, 12'd771, 12'd796, 12'd822, 12'd848, 12'd874, 12'd900, 12'd925, 12'd951, 12'd977, 12'd1003, 12'd1029, 12'd1054, 12'd1080, 12'd1106, 12'd1132, 12'd1158, 12'd1183, 12'd1209, 12'd1235, 12'd1261, 12'd1287, 12'd1312, 12'd1338, 12'd1364, 12'd1390, 12'd1416, 12'd1441, 12'd1467, 12'd1493, 12'd1519, 12'd1544, 12'd1570, 12'd1596, 12'd1622, 12'd1648, 12'd1673, 12'd1699, 12'd1725, 12'd1751, 12'd1777, 12'd1802, 12'd1828, 12'd1854, 12'd1880, 12'd1906, 12'd1931, 12'd1957, 12'd1983, 12'd2009, 12'd2035, 12'd2060, 12'd2086, 12'd2112, 12'd2138, 12'd2164, 12'd2189, 12'd2215, 12'd2241, 12'd2267, 12'd2293, 12'd2318, 12'd2344, 12'd2370, 12'd2396, 12'd2422, 12'd2447, 12'd2473, 12'd2499, 12'd2525, 12'd2551, 12'd2576, 12'd2602, 12'd2628, 12'd2654, 12'd2679, 12'd2705, 12'd2731, 12'd2757, 12'd2783, 12'd2808, 12'd2834, 12'd2860, 12'd2886, 12'd2912, 12'd2937, 12'd2963, 12'd2989, 12'd3015, 12'd3041, 12'd3066, 12'd3092, 12'd3118, 12'd3144, 12'd3170, 12'd3195, 12'd3221, 12'd3247, 12'd3273, 12'd3299, 12'd3324, 12'd3350, 12'd3376, 12'd3402, 12'd3428, 12'd3453, 12'd3479, 12'd3505, 12'd3531, 12'd3557, 12'd3582, 12'd3608, 12'd3634, 12'd3660, 12'd3686, 12'd3686, 12'd3660, 12'd3634, 12'd3608, 12'd3582, 12'd3557, 12'd3531, 12'd3505, 12'd3479, 12'd3453, 12'd3428, 12'd3402, 12'd3376, 12'd3350, 12'd3324, 12'd3299, 12'd3273, 12'd3247, 12'd3221, 12'd3195, 12'd3170, 12'd3144, 12'd3118, 12'd3092, 12'd3066, 12'd3041, 12'd3015, 12'd2989, 12'd2963, 12'd2937, 12'd2912, 12'd2886, 12'd2860, 12'd2834, 12'd2808, 12'd2783, 12'd2757, 12'd2731, 12'd2705, 12'd2679, 12'd2654, 12'd2628, 12'd2602, 12'd2576, 12'd2551, 12'd2525, 12'd2499, 12'd2473, 12'd2447, 12'd2422, 12'd2396, 12'd2370, 12'd2344, 12'd2318, 12'd2293, 12'd2267, 12'd2241, 12'd2215, 12'd2189, 12'd2164, 12'd2138, 12'd2112, 12'd2086, 12'd2060, 12'd2035, 12'd2009, 12'd1983, 12'd1957, 12'd1931, 12'd1906, 12'd1880, 12'd1854, 12'd1828, 12'd1802, 12'd1777, 12'd1751, 12'd1725, 12'd1699, 12'd1673, 12'd1648, 12'd1622, 12'd1596, 12'd1570, 12'd1544, 12'd1519, 12'd1493, 12'd1467, 12'd1441, 12'd1416, 12'd1390, 12'd1364, 12'd1338, 12'd1312, 12'd1287, 12'd1261, 12'd1235, 12'd1209, 12'd1183, 12'd1158, 12'd1132, 12'd1106, 12'd1080, 12'd1054, 12'd1029, 12'd1003, 12'd977, 12'd951, 12'd925, 12'd900, 12'd874, 12'd848, 12'd822, 12'd796, 12'd771, 12'd745, 12'd719, 12'd693, 12'd667, 12'd642, 12'd616, 12'd590, 12'd564, 12'd538, 12'd513, 12'd487, 12'd461, 12'd435, 12'd410 } ;
			// shape: triangle // depth: 5 //
			{ 3'd2, 3'd4 } : dataTable = { 12'd0, 12'd32, 12'd64, 12'd97, 12'd129, 12'd161, 12'd193, 12'd226, 12'd258, 12'd290, 12'd322, 12'd355, 12'd387, 12'd419, 12'd451, 12'd484, 12'd516, 12'd548, 12'd580, 12'd613, 12'd645, 12'd677, 12'd709, 12'd742, 12'd774, 12'd806, 12'd838, 12'd871, 12'd903, 12'd935, 12'd967, 12'd1000, 12'd1032, 12'd1064, 12'd1096, 12'd1129, 12'd1161, 12'd1193, 12'd1225, 12'd1258, 12'd1290, 12'd1322, 12'd1354, 12'd1386, 12'd1419, 12'd1451, 12'd1483, 12'd1515, 12'd1548, 12'd1580, 12'd1612, 12'd1644, 12'd1677, 12'd1709, 12'd1741, 12'd1773, 12'd1806, 12'd1838, 12'd1870, 12'd1902, 12'd1935, 12'd1967, 12'd1999, 12'd2031, 12'd2064, 12'd2096, 12'd2128, 12'd2160, 12'd2193, 12'd2225, 12'd2257, 12'd2289, 12'd2322, 12'd2354, 12'd2386, 12'd2418, 12'd2451, 12'd2483, 12'd2515, 12'd2547, 12'd2580, 12'd2612, 12'd2644, 12'd2676, 12'd2709, 12'd2741, 12'd2773, 12'd2805, 12'd2837, 12'd2870, 12'd2902, 12'd2934, 12'd2966, 12'd2999, 12'd3031, 12'd3063, 12'd3095, 12'd3128, 12'd3160, 12'd3192, 12'd3224, 12'd3257, 12'd3289, 12'd3321, 12'd3353, 12'd3386, 12'd3418, 12'd3450, 12'd3482, 12'd3515, 12'd3547, 12'd3579, 12'd3611, 12'd3644, 12'd3676, 12'd3708, 12'd3740, 12'd3773, 12'd3805, 12'd3837, 12'd3869, 12'd3902, 12'd3934, 12'd3966, 12'd3998, 12'd4031, 12'd4063, 12'd4095, 12'd4095, 12'd4063, 12'd4031, 12'd3998, 12'd3966, 12'd3934, 12'd3902, 12'd3869, 12'd3837, 12'd3805, 12'd3773, 12'd3740, 12'd3708, 12'd3676, 12'd3644, 12'd3611, 12'd3579, 12'd3547, 12'd3515, 12'd3482, 12'd3450, 12'd3418, 12'd3386, 12'd3353, 12'd3321, 12'd3289, 12'd3257, 12'd3224, 12'd3192, 12'd3160, 12'd3128, 12'd3095, 12'd3063, 12'd3031, 12'd2999, 12'd2966, 12'd2934, 12'd2902, 12'd2870, 12'd2837, 12'd2805, 12'd2773, 12'd2741, 12'd2709, 12'd2676, 12'd2644, 12'd2612, 12'd2580, 12'd2547, 12'd2515, 12'd2483, 12'd2451, 12'd2418, 12'd2386, 12'd2354, 12'd2322, 12'd2289, 12'd2257, 12'd2225, 12'd2193, 12'd2160, 12'd2128, 12'd2096, 12'd2064, 12'd2031, 12'd1999, 12'd1967, 12'd1935, 12'd1902, 12'd1870, 12'd1838, 12'd1806, 12'd1773, 12'd1741, 12'd1709, 12'd1677, 12'd1644, 12'd1612, 12'd1580, 12'd1548, 12'd1515, 12'd1483, 12'd1451, 12'd1419, 12'd1386, 12'd1354, 12'd1322, 12'd1290, 12'd1258, 12'd1225, 12'd1193, 12'd1161, 12'd1129, 12'd1096, 12'd1064, 12'd1032, 12'd1000, 12'd967, 12'd935, 12'd903, 12'd871, 12'd838, 12'd806, 12'd774, 12'd742, 12'd709, 12'd677, 12'd645, 12'd613, 12'd580, 12'd548, 12'd516, 12'd484, 12'd451, 12'd419, 12'd387, 12'd355, 12'd322, 12'd290, 12'd258, 12'd226, 12'd193, 12'd161, 12'd129, 12'd97, 12'd64, 12'd32, 12'd0 } ;
			// shape: ramp up // depth: 1 //
			{ 3'd3, 3'd0 } : dataTable = { 12'd1638, 12'd1641, 12'd1644, 12'd1648, 12'd1651, 12'd1654, 12'd1657, 12'd1660, 12'd1664, 12'd1667, 12'd1670, 12'd1673, 12'd1677, 12'd1680, 12'd1683, 12'd1686, 12'd1689, 12'd1693, 12'd1696, 12'd1699, 12'd1702, 12'd1705, 12'd1709, 12'd1712, 12'd1715, 12'd1718, 12'd1722, 12'd1725, 12'd1728, 12'd1731, 12'd1734, 12'd1738, 12'd1741, 12'd1744, 12'd1747, 12'd1750, 12'd1754, 12'd1757, 12'd1760, 12'd1763, 12'd1766, 12'd1770, 12'd1773, 12'd1776, 12'd1779, 12'd1783, 12'd1786, 12'd1789, 12'd1792, 12'd1795, 12'd1799, 12'd1802, 12'd1805, 12'd1808, 12'd1811, 12'd1815, 12'd1818, 12'd1821, 12'd1824, 12'd1827, 12'd1831, 12'd1834, 12'd1837, 12'd1840, 12'd1844, 12'd1847, 12'd1850, 12'd1853, 12'd1856, 12'd1860, 12'd1863, 12'd1866, 12'd1869, 12'd1872, 12'd1876, 12'd1879, 12'd1882, 12'd1885, 12'd1889, 12'd1892, 12'd1895, 12'd1898, 12'd1901, 12'd1905, 12'd1908, 12'd1911, 12'd1914, 12'd1917, 12'd1921, 12'd1924, 12'd1927, 12'd1930, 12'd1933, 12'd1937, 12'd1940, 12'd1943, 12'd1946, 12'd1950, 12'd1953, 12'd1956, 12'd1959, 12'd1962, 12'd1966, 12'd1969, 12'd1972, 12'd1975, 12'd1978, 12'd1982, 12'd1985, 12'd1988, 12'd1991, 12'd1995, 12'd1998, 12'd2001, 12'd2004, 12'd2007, 12'd2011, 12'd2014, 12'd2017, 12'd2020, 12'd2023, 12'd2027, 12'd2030, 12'd2033, 12'd2036, 12'd2039, 12'd2043, 12'd2046, 12'd2049, 12'd2052, 12'd2056, 12'd2059, 12'd2062, 12'd2065, 12'd2068, 12'd2072, 12'd2075, 12'd2078, 12'd2081, 12'd2084, 12'd2088, 12'd2091, 12'd2094, 12'd2097, 12'd2100, 12'd2104, 12'd2107, 12'd2110, 12'd2113, 12'd2117, 12'd2120, 12'd2123, 12'd2126, 12'd2129, 12'd2133, 12'd2136, 12'd2139, 12'd2142, 12'd2145, 12'd2149, 12'd2152, 12'd2155, 12'd2158, 12'd2162, 12'd2165, 12'd2168, 12'd2171, 12'd2174, 12'd2178, 12'd2181, 12'd2184, 12'd2187, 12'd2190, 12'd2194, 12'd2197, 12'd2200, 12'd2203, 12'd2206, 12'd2210, 12'd2213, 12'd2216, 12'd2219, 12'd2223, 12'd2226, 12'd2229, 12'd2232, 12'd2235, 12'd2239, 12'd2242, 12'd2245, 12'd2248, 12'd2251, 12'd2255, 12'd2258, 12'd2261, 12'd2264, 12'd2268, 12'd2271, 12'd2274, 12'd2277, 12'd2280, 12'd2284, 12'd2287, 12'd2290, 12'd2293, 12'd2296, 12'd2300, 12'd2303, 12'd2306, 12'd2309, 12'd2312, 12'd2316, 12'd2319, 12'd2322, 12'd2325, 12'd2329, 12'd2332, 12'd2335, 12'd2338, 12'd2341, 12'd2345, 12'd2348, 12'd2351, 12'd2354, 12'd2357, 12'd2361, 12'd2364, 12'd2367, 12'd2370, 12'd2373, 12'd2377, 12'd2380, 12'd2383, 12'd2386, 12'd2390, 12'd2393, 12'd2396, 12'd2399, 12'd2402, 12'd2406, 12'd2409, 12'd2412, 12'd2415, 12'd2418, 12'd2422, 12'd2425, 12'd2428, 12'd2431, 12'd2435, 12'd2438, 12'd2441, 12'd2444, 12'd2447, 12'd2451, 12'd2454, 12'd2457 } ;
			// shape: ramp up // depth: 2 //
			{ 3'd3, 3'd1 } : dataTable = { 12'd1228, 12'd1235, 12'd1241, 12'd1248, 12'd1254, 12'd1261, 12'd1267, 12'd1273, 12'd1280, 12'd1286, 12'd1293, 12'd1299, 12'd1306, 12'd1312, 12'd1318, 12'd1325, 12'd1331, 12'd1338, 12'd1344, 12'd1351, 12'd1357, 12'd1363, 12'd1370, 12'd1376, 12'd1383, 12'd1389, 12'd1396, 12'd1402, 12'd1408, 12'd1415, 12'd1421, 12'd1428, 12'd1434, 12'd1440, 12'd1447, 12'd1453, 12'd1460, 12'd1466, 12'd1473, 12'd1479, 12'd1485, 12'd1492, 12'd1498, 12'd1505, 12'd1511, 12'd1518, 12'd1524, 12'd1530, 12'd1537, 12'd1543, 12'd1550, 12'd1556, 12'd1563, 12'd1569, 12'd1575, 12'd1582, 12'd1588, 12'd1595, 12'd1601, 12'd1607, 12'd1614, 12'd1620, 12'd1627, 12'd1633, 12'd1640, 12'd1646, 12'd1652, 12'd1659, 12'd1665, 12'd1672, 12'd1678, 12'd1685, 12'd1691, 12'd1697, 12'd1704, 12'd1710, 12'd1717, 12'd1723, 12'd1730, 12'd1736, 12'd1742, 12'd1749, 12'd1755, 12'd1762, 12'd1768, 12'd1774, 12'd1781, 12'd1787, 12'd1794, 12'd1800, 12'd1807, 12'd1813, 12'd1819, 12'd1826, 12'd1832, 12'd1839, 12'd1845, 12'd1852, 12'd1858, 12'd1864, 12'd1871, 12'd1877, 12'd1884, 12'd1890, 12'd1897, 12'd1903, 12'd1909, 12'd1916, 12'd1922, 12'd1929, 12'd1935, 12'd1942, 12'd1948, 12'd1954, 12'd1961, 12'd1967, 12'd1974, 12'd1980, 12'd1986, 12'd1993, 12'd1999, 12'd2006, 12'd2012, 12'd2019, 12'd2025, 12'd2031, 12'd2038, 12'd2044, 12'd2051, 12'd2057, 12'd2064, 12'd2070, 12'd2076, 12'd2083, 12'd2089, 12'd2096, 12'd2102, 12'd2109, 12'd2115, 12'd2121, 12'd2128, 12'd2134, 12'd2141, 12'd2147, 12'd2153, 12'd2160, 12'd2166, 12'd2173, 12'd2179, 12'd2186, 12'd2192, 12'd2198, 12'd2205, 12'd2211, 12'd2218, 12'd2224, 12'd2231, 12'd2237, 12'd2243, 12'd2250, 12'd2256, 12'd2263, 12'd2269, 12'd2276, 12'd2282, 12'd2288, 12'd2295, 12'd2301, 12'd2308, 12'd2314, 12'd2320, 12'd2327, 12'd2333, 12'd2340, 12'd2346, 12'd2353, 12'd2359, 12'd2365, 12'd2372, 12'd2378, 12'd2385, 12'd2391, 12'd2398, 12'd2404, 12'd2410, 12'd2417, 12'd2423, 12'd2430, 12'd2436, 12'd2443, 12'd2449, 12'd2455, 12'd2462, 12'd2468, 12'd2475, 12'd2481, 12'd2488, 12'd2494, 12'd2500, 12'd2507, 12'd2513, 12'd2520, 12'd2526, 12'd2532, 12'd2539, 12'd2545, 12'd2552, 12'd2558, 12'd2565, 12'd2571, 12'd2577, 12'd2584, 12'd2590, 12'd2597, 12'd2603, 12'd2610, 12'd2616, 12'd2622, 12'd2629, 12'd2635, 12'd2642, 12'd2648, 12'd2655, 12'd2661, 12'd2667, 12'd2674, 12'd2680, 12'd2687, 12'd2693, 12'd2699, 12'd2706, 12'd2712, 12'd2719, 12'd2725, 12'd2732, 12'd2738, 12'd2744, 12'd2751, 12'd2757, 12'd2764, 12'd2770, 12'd2777, 12'd2783, 12'd2789, 12'd2796, 12'd2802, 12'd2809, 12'd2815, 12'd2822, 12'd2828, 12'd2834, 12'd2841, 12'd2847, 12'd2854, 12'd2860, 12'd2866 } ;
			// shape: ramp up // depth: 3 //
			{ 3'd3, 3'd2 } : dataTable = { 12'd819, 12'd829, 12'd838, 12'd848, 12'd858, 12'd867, 12'd877, 12'd886, 12'd896, 12'd906, 12'd915, 12'd925, 12'd935, 12'd944, 12'd954, 12'd964, 12'd973, 12'd983, 12'd992, 12'd1002, 12'd1012, 12'd1021, 12'd1031, 12'd1041, 12'd1050, 12'd1060, 12'd1070, 12'd1079, 12'd1089, 12'd1098, 12'd1108, 12'd1118, 12'd1127, 12'd1137, 12'd1147, 12'd1156, 12'd1166, 12'd1176, 12'd1185, 12'd1195, 12'd1204, 12'd1214, 12'd1224, 12'd1233, 12'd1243, 12'd1253, 12'd1262, 12'd1272, 12'd1281, 12'd1291, 12'd1301, 12'd1310, 12'd1320, 12'd1330, 12'd1339, 12'd1349, 12'd1359, 12'd1368, 12'd1378, 12'd1387, 12'd1397, 12'd1407, 12'd1416, 12'd1426, 12'd1436, 12'd1445, 12'd1455, 12'd1465, 12'd1474, 12'd1484, 12'd1493, 12'd1503, 12'd1513, 12'd1522, 12'd1532, 12'd1542, 12'd1551, 12'd1561, 12'd1571, 12'd1580, 12'd1590, 12'd1599, 12'd1609, 12'd1619, 12'd1628, 12'd1638, 12'd1648, 12'd1657, 12'd1667, 12'd1677, 12'd1686, 12'd1696, 12'd1705, 12'd1715, 12'd1725, 12'd1734, 12'd1744, 12'd1754, 12'd1763, 12'd1773, 12'd1783, 12'd1792, 12'd1802, 12'd1811, 12'd1821, 12'd1831, 12'd1840, 12'd1850, 12'd1860, 12'd1869, 12'd1879, 12'd1889, 12'd1898, 12'd1908, 12'd1917, 12'd1927, 12'd1937, 12'd1946, 12'd1956, 12'd1966, 12'd1975, 12'd1985, 12'd1995, 12'd2004, 12'd2014, 12'd2023, 12'd2033, 12'd2043, 12'd2052, 12'd2062, 12'd2072, 12'd2081, 12'd2091, 12'd2100, 12'd2110, 12'd2120, 12'd2129, 12'd2139, 12'd2149, 12'd2158, 12'd2168, 12'd2178, 12'd2187, 12'd2197, 12'd2206, 12'd2216, 12'd2226, 12'd2235, 12'd2245, 12'd2255, 12'd2264, 12'd2274, 12'd2284, 12'd2293, 12'd2303, 12'd2312, 12'd2322, 12'd2332, 12'd2341, 12'd2351, 12'd2361, 12'd2370, 12'd2380, 12'd2390, 12'd2399, 12'd2409, 12'd2418, 12'd2428, 12'd2438, 12'd2447, 12'd2457, 12'd2467, 12'd2476, 12'd2486, 12'd2496, 12'd2505, 12'd2515, 12'd2524, 12'd2534, 12'd2544, 12'd2553, 12'd2563, 12'd2573, 12'd2582, 12'd2592, 12'd2602, 12'd2611, 12'd2621, 12'd2630, 12'd2640, 12'd2650, 12'd2659, 12'd2669, 12'd2679, 12'd2688, 12'd2698, 12'd2708, 12'd2717, 12'd2727, 12'd2736, 12'd2746, 12'd2756, 12'd2765, 12'd2775, 12'd2785, 12'd2794, 12'd2804, 12'd2814, 12'd2823, 12'd2833, 12'd2842, 12'd2852, 12'd2862, 12'd2871, 12'd2881, 12'd2891, 12'd2900, 12'd2910, 12'd2919, 12'd2929, 12'd2939, 12'd2948, 12'd2958, 12'd2968, 12'd2977, 12'd2987, 12'd2997, 12'd3006, 12'd3016, 12'd3025, 12'd3035, 12'd3045, 12'd3054, 12'd3064, 12'd3074, 12'd3083, 12'd3093, 12'd3103, 12'd3112, 12'd3122, 12'd3131, 12'd3141, 12'd3151, 12'd3160, 12'd3170, 12'd3180, 12'd3189, 12'd3199, 12'd3209, 12'd3218, 12'd3228, 12'd3237, 12'd3247, 12'd3257, 12'd3266, 12'd3276 } ;
			// shape: ramp up // depth: 4 //
			{ 3'd3, 3'd3 } : dataTable = { 12'd410, 12'd422, 12'd435, 12'd448, 12'd461, 12'd474, 12'd487, 12'd499, 12'd512, 12'd525, 12'd538, 12'd551, 12'd564, 12'd577, 12'd589, 12'd602, 12'd615, 12'd628, 12'd641, 12'd654, 12'd666, 12'd679, 12'd692, 12'd705, 12'd718, 12'd731, 12'd744, 12'd756, 12'd769, 12'd782, 12'd795, 12'd808, 12'd821, 12'd833, 12'd846, 12'd859, 12'd872, 12'd885, 12'd898, 12'd911, 12'd923, 12'd936, 12'd949, 12'd962, 12'd975, 12'd988, 12'd1000, 12'd1013, 12'd1026, 12'd1039, 12'd1052, 12'd1065, 12'd1078, 12'd1090, 12'd1103, 12'd1116, 12'd1129, 12'd1142, 12'd1155, 12'd1167, 12'd1180, 12'd1193, 12'd1206, 12'd1219, 12'd1232, 12'd1245, 12'd1257, 12'd1270, 12'd1283, 12'd1296, 12'd1309, 12'd1322, 12'd1334, 12'd1347, 12'd1360, 12'd1373, 12'd1386, 12'd1399, 12'd1412, 12'd1424, 12'd1437, 12'd1450, 12'd1463, 12'd1476, 12'd1489, 12'd1502, 12'd1514, 12'd1527, 12'd1540, 12'd1553, 12'd1566, 12'd1579, 12'd1591, 12'd1604, 12'd1617, 12'd1630, 12'd1643, 12'd1656, 12'd1669, 12'd1681, 12'd1694, 12'd1707, 12'd1720, 12'd1733, 12'd1746, 12'd1758, 12'd1771, 12'd1784, 12'd1797, 12'd1810, 12'd1823, 12'd1836, 12'd1848, 12'd1861, 12'd1874, 12'd1887, 12'd1900, 12'd1913, 12'd1925, 12'd1938, 12'd1951, 12'd1964, 12'd1977, 12'd1990, 12'd2003, 12'd2015, 12'd2028, 12'd2041, 12'd2054, 12'd2067, 12'd2080, 12'd2092, 12'd2105, 12'd2118, 12'd2131, 12'd2144, 12'd2157, 12'd2170, 12'd2182, 12'd2195, 12'd2208, 12'd2221, 12'd2234, 12'd2247, 12'd2259, 12'd2272, 12'd2285, 12'd2298, 12'd2311, 12'd2324, 12'd2337, 12'd2349, 12'd2362, 12'd2375, 12'd2388, 12'd2401, 12'd2414, 12'd2426, 12'd2439, 12'd2452, 12'd2465, 12'd2478, 12'd2491, 12'd2504, 12'd2516, 12'd2529, 12'd2542, 12'd2555, 12'd2568, 12'd2581, 12'd2594, 12'd2606, 12'd2619, 12'd2632, 12'd2645, 12'd2658, 12'd2671, 12'd2683, 12'd2696, 12'd2709, 12'd2722, 12'd2735, 12'd2748, 12'd2761, 12'd2773, 12'd2786, 12'd2799, 12'd2812, 12'd2825, 12'd2838, 12'd2850, 12'd2863, 12'd2876, 12'd2889, 12'd2902, 12'd2915, 12'd2928, 12'd2940, 12'd2953, 12'd2966, 12'd2979, 12'd2992, 12'd3005, 12'd3017, 12'd3030, 12'd3043, 12'd3056, 12'd3069, 12'd3082, 12'd3095, 12'd3107, 12'd3120, 12'd3133, 12'd3146, 12'd3159, 12'd3172, 12'd3184, 12'd3197, 12'd3210, 12'd3223, 12'd3236, 12'd3249, 12'd3262, 12'd3274, 12'd3287, 12'd3300, 12'd3313, 12'd3326, 12'd3339, 12'd3351, 12'd3364, 12'd3377, 12'd3390, 12'd3403, 12'd3416, 12'd3429, 12'd3441, 12'd3454, 12'd3467, 12'd3480, 12'd3493, 12'd3506, 12'd3518, 12'd3531, 12'd3544, 12'd3557, 12'd3570, 12'd3583, 12'd3596, 12'd3608, 12'd3621, 12'd3634, 12'd3647, 12'd3660, 12'd3673, 12'd3686 } ;
			// shape: ramp up // depth: 5 //
			{ 3'd3, 3'd4 } : dataTable = { 12'd0, 12'd16, 12'd32, 12'd48, 12'd64, 12'd80, 12'd96, 12'd112, 12'd128, 12'd145, 12'd161, 12'd177, 12'd193, 12'd209, 12'd225, 12'd241, 12'd257, 12'd273, 12'd289, 12'd305, 12'd321, 12'd337, 12'd353, 12'd369, 12'd385, 12'd401, 12'd418, 12'd434, 12'd450, 12'd466, 12'd482, 12'd498, 12'd514, 12'd530, 12'd546, 12'd562, 12'd578, 12'd594, 12'd610, 12'd626, 12'd642, 12'd658, 12'd674, 12'd691, 12'd707, 12'd723, 12'd739, 12'd755, 12'd771, 12'd787, 12'd803, 12'd819, 12'd835, 12'd851, 12'd867, 12'd883, 12'd899, 12'd915, 12'd931, 12'd947, 12'd964, 12'd980, 12'd996, 12'd1012, 12'd1028, 12'd1044, 12'd1060, 12'd1076, 12'd1092, 12'd1108, 12'd1124, 12'd1140, 12'd1156, 12'd1172, 12'd1188, 12'd1204, 12'd1220, 12'd1237, 12'd1253, 12'd1269, 12'd1285, 12'd1301, 12'd1317, 12'd1333, 12'd1349, 12'd1365, 12'd1381, 12'd1397, 12'd1413, 12'd1429, 12'd1445, 12'd1461, 12'd1477, 12'd1493, 12'd1510, 12'd1526, 12'd1542, 12'd1558, 12'd1574, 12'd1590, 12'd1606, 12'd1622, 12'd1638, 12'd1654, 12'd1670, 12'd1686, 12'd1702, 12'd1718, 12'd1734, 12'd1750, 12'd1766, 12'd1783, 12'd1799, 12'd1815, 12'd1831, 12'd1847, 12'd1863, 12'd1879, 12'd1895, 12'd1911, 12'd1927, 12'd1943, 12'd1959, 12'd1975, 12'd1991, 12'd2007, 12'd2023, 12'd2039, 12'd2056, 12'd2072, 12'd2088, 12'd2104, 12'd2120, 12'd2136, 12'd2152, 12'd2168, 12'd2184, 12'd2200, 12'd2216, 12'd2232, 12'd2248, 12'd2264, 12'd2280, 12'd2296, 12'd2312, 12'd2329, 12'd2345, 12'd2361, 12'd2377, 12'd2393, 12'd2409, 12'd2425, 12'd2441, 12'd2457, 12'd2473, 12'd2489, 12'd2505, 12'd2521, 12'd2537, 12'd2553, 12'd2569, 12'd2585, 12'd2602, 12'd2618, 12'd2634, 12'd2650, 12'd2666, 12'd2682, 12'd2698, 12'd2714, 12'd2730, 12'd2746, 12'd2762, 12'd2778, 12'd2794, 12'd2810, 12'd2826, 12'd2842, 12'd2858, 12'd2875, 12'd2891, 12'd2907, 12'd2923, 12'd2939, 12'd2955, 12'd2971, 12'd2987, 12'd3003, 12'd3019, 12'd3035, 12'd3051, 12'd3067, 12'd3083, 12'd3099, 12'd3115, 12'd3131, 12'd3148, 12'd3164, 12'd3180, 12'd3196, 12'd3212, 12'd3228, 12'd3244, 12'd3260, 12'd3276, 12'd3292, 12'd3308, 12'd3324, 12'd3340, 12'd3356, 12'd3372, 12'd3388, 12'd3404, 12'd3421, 12'd3437, 12'd3453, 12'd3469, 12'd3485, 12'd3501, 12'd3517, 12'd3533, 12'd3549, 12'd3565, 12'd3581, 12'd3597, 12'd3613, 12'd3629, 12'd3645, 12'd3661, 12'd3677, 12'd3694, 12'd3710, 12'd3726, 12'd3742, 12'd3758, 12'd3774, 12'd3790, 12'd3806, 12'd3822, 12'd3838, 12'd3854, 12'd3870, 12'd3886, 12'd3902, 12'd3918, 12'd3934, 12'd3950, 12'd3967, 12'd3983, 12'd3999, 12'd4015, 12'd4031, 12'd4047, 12'd4063, 12'd4079, 12'd4095 } ;
			// shape: ramp down // depth: 1 //
			{ 3'd4, 3'd0 } : dataTable = { 12'd2457, 12'd2454, 12'd2451, 12'd2447, 12'd2444, 12'd2441, 12'd2438, 12'd2435, 12'd2431, 12'd2428, 12'd2425, 12'd2422, 12'd2418, 12'd2415, 12'd2412, 12'd2409, 12'd2406, 12'd2402, 12'd2399, 12'd2396, 12'd2393, 12'd2390, 12'd2386, 12'd2383, 12'd2380, 12'd2377, 12'd2373, 12'd2370, 12'd2367, 12'd2364, 12'd2361, 12'd2357, 12'd2354, 12'd2351, 12'd2348, 12'd2345, 12'd2341, 12'd2338, 12'd2335, 12'd2332, 12'd2329, 12'd2325, 12'd2322, 12'd2319, 12'd2316, 12'd2312, 12'd2309, 12'd2306, 12'd2303, 12'd2300, 12'd2296, 12'd2293, 12'd2290, 12'd2287, 12'd2284, 12'd2280, 12'd2277, 12'd2274, 12'd2271, 12'd2268, 12'd2264, 12'd2261, 12'd2258, 12'd2255, 12'd2251, 12'd2248, 12'd2245, 12'd2242, 12'd2239, 12'd2235, 12'd2232, 12'd2229, 12'd2226, 12'd2223, 12'd2219, 12'd2216, 12'd2213, 12'd2210, 12'd2206, 12'd2203, 12'd2200, 12'd2197, 12'd2194, 12'd2190, 12'd2187, 12'd2184, 12'd2181, 12'd2178, 12'd2174, 12'd2171, 12'd2168, 12'd2165, 12'd2162, 12'd2158, 12'd2155, 12'd2152, 12'd2149, 12'd2145, 12'd2142, 12'd2139, 12'd2136, 12'd2133, 12'd2129, 12'd2126, 12'd2123, 12'd2120, 12'd2117, 12'd2113, 12'd2110, 12'd2107, 12'd2104, 12'd2100, 12'd2097, 12'd2094, 12'd2091, 12'd2088, 12'd2084, 12'd2081, 12'd2078, 12'd2075, 12'd2072, 12'd2068, 12'd2065, 12'd2062, 12'd2059, 12'd2056, 12'd2052, 12'd2049, 12'd2046, 12'd2043, 12'd2039, 12'd2036, 12'd2033, 12'd2030, 12'd2027, 12'd2023, 12'd2020, 12'd2017, 12'd2014, 12'd2011, 12'd2007, 12'd2004, 12'd2001, 12'd1998, 12'd1995, 12'd1991, 12'd1988, 12'd1985, 12'd1982, 12'd1978, 12'd1975, 12'd1972, 12'd1969, 12'd1966, 12'd1962, 12'd1959, 12'd1956, 12'd1953, 12'd1950, 12'd1946, 12'd1943, 12'd1940, 12'd1937, 12'd1933, 12'd1930, 12'd1927, 12'd1924, 12'd1921, 12'd1917, 12'd1914, 12'd1911, 12'd1908, 12'd1905, 12'd1901, 12'd1898, 12'd1895, 12'd1892, 12'd1889, 12'd1885, 12'd1882, 12'd1879, 12'd1876, 12'd1872, 12'd1869, 12'd1866, 12'd1863, 12'd1860, 12'd1856, 12'd1853, 12'd1850, 12'd1847, 12'd1844, 12'd1840, 12'd1837, 12'd1834, 12'd1831, 12'd1827, 12'd1824, 12'd1821, 12'd1818, 12'd1815, 12'd1811, 12'd1808, 12'd1805, 12'd1802, 12'd1799, 12'd1795, 12'd1792, 12'd1789, 12'd1786, 12'd1783, 12'd1779, 12'd1776, 12'd1773, 12'd1770, 12'd1766, 12'd1763, 12'd1760, 12'd1757, 12'd1754, 12'd1750, 12'd1747, 12'd1744, 12'd1741, 12'd1738, 12'd1734, 12'd1731, 12'd1728, 12'd1725, 12'd1722, 12'd1718, 12'd1715, 12'd1712, 12'd1709, 12'd1705, 12'd1702, 12'd1699, 12'd1696, 12'd1693, 12'd1689, 12'd1686, 12'd1683, 12'd1680, 12'd1677, 12'd1673, 12'd1670, 12'd1667, 12'd1664, 12'd1660, 12'd1657, 12'd1654, 12'd1651, 12'd1648, 12'd1644, 12'd1641, 12'd1638 } ;
			// shape: ramp down // depth: 2 //
			{ 3'd4, 3'd1 } : dataTable = { 12'd2866, 12'd2860, 12'd2854, 12'd2847, 12'd2841, 12'd2834, 12'd2828, 12'd2822, 12'd2815, 12'd2809, 12'd2802, 12'd2796, 12'd2789, 12'd2783, 12'd2777, 12'd2770, 12'd2764, 12'd2757, 12'd2751, 12'd2744, 12'd2738, 12'd2732, 12'd2725, 12'd2719, 12'd2712, 12'd2706, 12'd2699, 12'd2693, 12'd2687, 12'd2680, 12'd2674, 12'd2667, 12'd2661, 12'd2655, 12'd2648, 12'd2642, 12'd2635, 12'd2629, 12'd2622, 12'd2616, 12'd2610, 12'd2603, 12'd2597, 12'd2590, 12'd2584, 12'd2577, 12'd2571, 12'd2565, 12'd2558, 12'd2552, 12'd2545, 12'd2539, 12'd2532, 12'd2526, 12'd2520, 12'd2513, 12'd2507, 12'd2500, 12'd2494, 12'd2488, 12'd2481, 12'd2475, 12'd2468, 12'd2462, 12'd2455, 12'd2449, 12'd2443, 12'd2436, 12'd2430, 12'd2423, 12'd2417, 12'd2410, 12'd2404, 12'd2398, 12'd2391, 12'd2385, 12'd2378, 12'd2372, 12'd2365, 12'd2359, 12'd2353, 12'd2346, 12'd2340, 12'd2333, 12'd2327, 12'd2320, 12'd2314, 12'd2308, 12'd2301, 12'd2295, 12'd2288, 12'd2282, 12'd2276, 12'd2269, 12'd2263, 12'd2256, 12'd2250, 12'd2243, 12'd2237, 12'd2231, 12'd2224, 12'd2218, 12'd2211, 12'd2205, 12'd2198, 12'd2192, 12'd2186, 12'd2179, 12'd2173, 12'd2166, 12'd2160, 12'd2153, 12'd2147, 12'd2141, 12'd2134, 12'd2128, 12'd2121, 12'd2115, 12'd2109, 12'd2102, 12'd2096, 12'd2089, 12'd2083, 12'd2076, 12'd2070, 12'd2064, 12'd2057, 12'd2051, 12'd2044, 12'd2038, 12'd2031, 12'd2025, 12'd2019, 12'd2012, 12'd2006, 12'd1999, 12'd1993, 12'd1986, 12'd1980, 12'd1974, 12'd1967, 12'd1961, 12'd1954, 12'd1948, 12'd1942, 12'd1935, 12'd1929, 12'd1922, 12'd1916, 12'd1909, 12'd1903, 12'd1897, 12'd1890, 12'd1884, 12'd1877, 12'd1871, 12'd1864, 12'd1858, 12'd1852, 12'd1845, 12'd1839, 12'd1832, 12'd1826, 12'd1819, 12'd1813, 12'd1807, 12'd1800, 12'd1794, 12'd1787, 12'd1781, 12'd1775, 12'd1768, 12'd1762, 12'd1755, 12'd1749, 12'd1742, 12'd1736, 12'd1730, 12'd1723, 12'd1717, 12'd1710, 12'd1704, 12'd1697, 12'd1691, 12'd1685, 12'd1678, 12'd1672, 12'd1665, 12'd1659, 12'd1652, 12'd1646, 12'd1640, 12'd1633, 12'd1627, 12'd1620, 12'd1614, 12'd1607, 12'd1601, 12'd1595, 12'd1588, 12'd1582, 12'd1575, 12'd1569, 12'd1563, 12'd1556, 12'd1550, 12'd1543, 12'd1537, 12'd1530, 12'd1524, 12'd1518, 12'd1511, 12'd1505, 12'd1498, 12'd1492, 12'd1485, 12'd1479, 12'd1473, 12'd1466, 12'd1460, 12'd1453, 12'd1447, 12'd1440, 12'd1434, 12'd1428, 12'd1421, 12'd1415, 12'd1408, 12'd1402, 12'd1396, 12'd1389, 12'd1383, 12'd1376, 12'd1370, 12'd1363, 12'd1357, 12'd1351, 12'd1344, 12'd1338, 12'd1331, 12'd1325, 12'd1318, 12'd1312, 12'd1306, 12'd1299, 12'd1293, 12'd1286, 12'd1280, 12'd1273, 12'd1267, 12'd1261, 12'd1254, 12'd1248, 12'd1241, 12'd1235, 12'd1228 } ;
			// shape: ramp down // depth: 3 //
			{ 3'd4, 3'd2 } : dataTable = { 12'd3276, 12'd3266, 12'd3257, 12'd3247, 12'd3237, 12'd3228, 12'd3218, 12'd3209, 12'd3199, 12'd3189, 12'd3180, 12'd3170, 12'd3160, 12'd3151, 12'd3141, 12'd3131, 12'd3122, 12'd3112, 12'd3103, 12'd3093, 12'd3083, 12'd3074, 12'd3064, 12'd3054, 12'd3045, 12'd3035, 12'd3025, 12'd3016, 12'd3006, 12'd2997, 12'd2987, 12'd2977, 12'd2968, 12'd2958, 12'd2948, 12'd2939, 12'd2929, 12'd2919, 12'd2910, 12'd2900, 12'd2891, 12'd2881, 12'd2871, 12'd2862, 12'd2852, 12'd2842, 12'd2833, 12'd2823, 12'd2814, 12'd2804, 12'd2794, 12'd2785, 12'd2775, 12'd2765, 12'd2756, 12'd2746, 12'd2736, 12'd2727, 12'd2717, 12'd2708, 12'd2698, 12'd2688, 12'd2679, 12'd2669, 12'd2659, 12'd2650, 12'd2640, 12'd2630, 12'd2621, 12'd2611, 12'd2602, 12'd2592, 12'd2582, 12'd2573, 12'd2563, 12'd2553, 12'd2544, 12'd2534, 12'd2524, 12'd2515, 12'd2505, 12'd2496, 12'd2486, 12'd2476, 12'd2467, 12'd2457, 12'd2447, 12'd2438, 12'd2428, 12'd2418, 12'd2409, 12'd2399, 12'd2390, 12'd2380, 12'd2370, 12'd2361, 12'd2351, 12'd2341, 12'd2332, 12'd2322, 12'd2312, 12'd2303, 12'd2293, 12'd2284, 12'd2274, 12'd2264, 12'd2255, 12'd2245, 12'd2235, 12'd2226, 12'd2216, 12'd2206, 12'd2197, 12'd2187, 12'd2178, 12'd2168, 12'd2158, 12'd2149, 12'd2139, 12'd2129, 12'd2120, 12'd2110, 12'd2100, 12'd2091, 12'd2081, 12'd2072, 12'd2062, 12'd2052, 12'd2043, 12'd2033, 12'd2023, 12'd2014, 12'd2004, 12'd1995, 12'd1985, 12'd1975, 12'd1966, 12'd1956, 12'd1946, 12'd1937, 12'd1927, 12'd1917, 12'd1908, 12'd1898, 12'd1889, 12'd1879, 12'd1869, 12'd1860, 12'd1850, 12'd1840, 12'd1831, 12'd1821, 12'd1811, 12'd1802, 12'd1792, 12'd1783, 12'd1773, 12'd1763, 12'd1754, 12'd1744, 12'd1734, 12'd1725, 12'd1715, 12'd1705, 12'd1696, 12'd1686, 12'd1677, 12'd1667, 12'd1657, 12'd1648, 12'd1638, 12'd1628, 12'd1619, 12'd1609, 12'd1599, 12'd1590, 12'd1580, 12'd1571, 12'd1561, 12'd1551, 12'd1542, 12'd1532, 12'd1522, 12'd1513, 12'd1503, 12'd1493, 12'd1484, 12'd1474, 12'd1465, 12'd1455, 12'd1445, 12'd1436, 12'd1426, 12'd1416, 12'd1407, 12'd1397, 12'd1387, 12'd1378, 12'd1368, 12'd1359, 12'd1349, 12'd1339, 12'd1330, 12'd1320, 12'd1310, 12'd1301, 12'd1291, 12'd1281, 12'd1272, 12'd1262, 12'd1253, 12'd1243, 12'd1233, 12'd1224, 12'd1214, 12'd1204, 12'd1195, 12'd1185, 12'd1176, 12'd1166, 12'd1156, 12'd1147, 12'd1137, 12'd1127, 12'd1118, 12'd1108, 12'd1098, 12'd1089, 12'd1079, 12'd1070, 12'd1060, 12'd1050, 12'd1041, 12'd1031, 12'd1021, 12'd1012, 12'd1002, 12'd992, 12'd983, 12'd973, 12'd964, 12'd954, 12'd944, 12'd935, 12'd925, 12'd915, 12'd906, 12'd896, 12'd886, 12'd877, 12'd867, 12'd858, 12'd848, 12'd838, 12'd829, 12'd819 } ;
			// shape: ramp down // depth: 4 //
			{ 3'd4, 3'd3 } : dataTable = { 12'd3686, 12'd3673, 12'd3660, 12'd3647, 12'd3634, 12'd3621, 12'd3608, 12'd3596, 12'd3583, 12'd3570, 12'd3557, 12'd3544, 12'd3531, 12'd3518, 12'd3506, 12'd3493, 12'd3480, 12'd3467, 12'd3454, 12'd3441, 12'd3429, 12'd3416, 12'd3403, 12'd3390, 12'd3377, 12'd3364, 12'd3351, 12'd3339, 12'd3326, 12'd3313, 12'd3300, 12'd3287, 12'd3274, 12'd3262, 12'd3249, 12'd3236, 12'd3223, 12'd3210, 12'd3197, 12'd3184, 12'd3172, 12'd3159, 12'd3146, 12'd3133, 12'd3120, 12'd3107, 12'd3095, 12'd3082, 12'd3069, 12'd3056, 12'd3043, 12'd3030, 12'd3017, 12'd3005, 12'd2992, 12'd2979, 12'd2966, 12'd2953, 12'd2940, 12'd2928, 12'd2915, 12'd2902, 12'd2889, 12'd2876, 12'd2863, 12'd2850, 12'd2838, 12'd2825, 12'd2812, 12'd2799, 12'd2786, 12'd2773, 12'd2761, 12'd2748, 12'd2735, 12'd2722, 12'd2709, 12'd2696, 12'd2683, 12'd2671, 12'd2658, 12'd2645, 12'd2632, 12'd2619, 12'd2606, 12'd2594, 12'd2581, 12'd2568, 12'd2555, 12'd2542, 12'd2529, 12'd2516, 12'd2504, 12'd2491, 12'd2478, 12'd2465, 12'd2452, 12'd2439, 12'd2426, 12'd2414, 12'd2401, 12'd2388, 12'd2375, 12'd2362, 12'd2349, 12'd2337, 12'd2324, 12'd2311, 12'd2298, 12'd2285, 12'd2272, 12'd2259, 12'd2247, 12'd2234, 12'd2221, 12'd2208, 12'd2195, 12'd2182, 12'd2170, 12'd2157, 12'd2144, 12'd2131, 12'd2118, 12'd2105, 12'd2092, 12'd2080, 12'd2067, 12'd2054, 12'd2041, 12'd2028, 12'd2015, 12'd2003, 12'd1990, 12'd1977, 12'd1964, 12'd1951, 12'd1938, 12'd1925, 12'd1913, 12'd1900, 12'd1887, 12'd1874, 12'd1861, 12'd1848, 12'd1836, 12'd1823, 12'd1810, 12'd1797, 12'd1784, 12'd1771, 12'd1758, 12'd1746, 12'd1733, 12'd1720, 12'd1707, 12'd1694, 12'd1681, 12'd1669, 12'd1656, 12'd1643, 12'd1630, 12'd1617, 12'd1604, 12'd1591, 12'd1579, 12'd1566, 12'd1553, 12'd1540, 12'd1527, 12'd1514, 12'd1502, 12'd1489, 12'd1476, 12'd1463, 12'd1450, 12'd1437, 12'd1424, 12'd1412, 12'd1399, 12'd1386, 12'd1373, 12'd1360, 12'd1347, 12'd1334, 12'd1322, 12'd1309, 12'd1296, 12'd1283, 12'd1270, 12'd1257, 12'd1245, 12'd1232, 12'd1219, 12'd1206, 12'd1193, 12'd1180, 12'd1167, 12'd1155, 12'd1142, 12'd1129, 12'd1116, 12'd1103, 12'd1090, 12'd1078, 12'd1065, 12'd1052, 12'd1039, 12'd1026, 12'd1013, 12'd1000, 12'd988, 12'd975, 12'd962, 12'd949, 12'd936, 12'd923, 12'd911, 12'd898, 12'd885, 12'd872, 12'd859, 12'd846, 12'd833, 12'd821, 12'd808, 12'd795, 12'd782, 12'd769, 12'd756, 12'd744, 12'd731, 12'd718, 12'd705, 12'd692, 12'd679, 12'd666, 12'd654, 12'd641, 12'd628, 12'd615, 12'd602, 12'd589, 12'd577, 12'd564, 12'd551, 12'd538, 12'd525, 12'd512, 12'd499, 12'd487, 12'd474, 12'd461, 12'd448, 12'd435, 12'd422, 12'd410 } ;
			// shape: ramp down // depth: 5 //
			{ 3'd4, 3'd4 } : dataTable = { 12'd4095, 12'd4079, 12'd4063, 12'd4047, 12'd4031, 12'd4015, 12'd3999, 12'd3983, 12'd3967, 12'd3950, 12'd3934, 12'd3918, 12'd3902, 12'd3886, 12'd3870, 12'd3854, 12'd3838, 12'd3822, 12'd3806, 12'd3790, 12'd3774, 12'd3758, 12'd3742, 12'd3726, 12'd3710, 12'd3694, 12'd3677, 12'd3661, 12'd3645, 12'd3629, 12'd3613, 12'd3597, 12'd3581, 12'd3565, 12'd3549, 12'd3533, 12'd3517, 12'd3501, 12'd3485, 12'd3469, 12'd3453, 12'd3437, 12'd3421, 12'd3404, 12'd3388, 12'd3372, 12'd3356, 12'd3340, 12'd3324, 12'd3308, 12'd3292, 12'd3276, 12'd3260, 12'd3244, 12'd3228, 12'd3212, 12'd3196, 12'd3180, 12'd3164, 12'd3148, 12'd3131, 12'd3115, 12'd3099, 12'd3083, 12'd3067, 12'd3051, 12'd3035, 12'd3019, 12'd3003, 12'd2987, 12'd2971, 12'd2955, 12'd2939, 12'd2923, 12'd2907, 12'd2891, 12'd2875, 12'd2858, 12'd2842, 12'd2826, 12'd2810, 12'd2794, 12'd2778, 12'd2762, 12'd2746, 12'd2730, 12'd2714, 12'd2698, 12'd2682, 12'd2666, 12'd2650, 12'd2634, 12'd2618, 12'd2602, 12'd2585, 12'd2569, 12'd2553, 12'd2537, 12'd2521, 12'd2505, 12'd2489, 12'd2473, 12'd2457, 12'd2441, 12'd2425, 12'd2409, 12'd2393, 12'd2377, 12'd2361, 12'd2345, 12'd2329, 12'd2312, 12'd2296, 12'd2280, 12'd2264, 12'd2248, 12'd2232, 12'd2216, 12'd2200, 12'd2184, 12'd2168, 12'd2152, 12'd2136, 12'd2120, 12'd2104, 12'd2088, 12'd2072, 12'd2056, 12'd2039, 12'd2023, 12'd2007, 12'd1991, 12'd1975, 12'd1959, 12'd1943, 12'd1927, 12'd1911, 12'd1895, 12'd1879, 12'd1863, 12'd1847, 12'd1831, 12'd1815, 12'd1799, 12'd1783, 12'd1766, 12'd1750, 12'd1734, 12'd1718, 12'd1702, 12'd1686, 12'd1670, 12'd1654, 12'd1638, 12'd1622, 12'd1606, 12'd1590, 12'd1574, 12'd1558, 12'd1542, 12'd1526, 12'd1510, 12'd1493, 12'd1477, 12'd1461, 12'd1445, 12'd1429, 12'd1413, 12'd1397, 12'd1381, 12'd1365, 12'd1349, 12'd1333, 12'd1317, 12'd1301, 12'd1285, 12'd1269, 12'd1253, 12'd1237, 12'd1220, 12'd1204, 12'd1188, 12'd1172, 12'd1156, 12'd1140, 12'd1124, 12'd1108, 12'd1092, 12'd1076, 12'd1060, 12'd1044, 12'd1028, 12'd1012, 12'd996, 12'd980, 12'd964, 12'd947, 12'd931, 12'd915, 12'd899, 12'd883, 12'd867, 12'd851, 12'd835, 12'd819, 12'd803, 12'd787, 12'd771, 12'd755, 12'd739, 12'd723, 12'd707, 12'd691, 12'd674, 12'd658, 12'd642, 12'd626, 12'd610, 12'd594, 12'd578, 12'd562, 12'd546, 12'd530, 12'd514, 12'd498, 12'd482, 12'd466, 12'd450, 12'd434, 12'd418, 12'd401, 12'd385, 12'd369, 12'd353, 12'd337, 12'd321, 12'd305, 12'd289, 12'd273, 12'd257, 12'd241, 12'd225, 12'd209, 12'd193, 12'd177, 12'd161, 12'd145, 12'd128, 12'd112, 12'd96, 12'd80, 12'd64, 12'd48, 12'd32, 12'd16, 12'd0 } ;
			default : dataTable = '0 ;
		endcase
	end

	// assign randomly generated index values for sample & hold
	assign SnH_index = { 8'd139, 8'd184, 8'd134, 8'd254, 8'd56, 8'd27, 8'd28, 8'd17, 8'd104, 8'd115, 8'd94, 8'd195, 8'd161, 8'd197, 8'd238, 8'd249, 8'd49, 8'd36, 8'd178, 8'd24, 8'd134, 8'd136, 8'd220, 8'd124, 8'd101, 8'd172, 8'd190, 8'd133, 8'd89, 8'd39, 8'd150, 8'd67, 8'd12, 8'd193, 8'd62, 8'd113, 8'd176, 8'd92, 8'd188, 8'd101, 8'd175, 8'd180, 8'd113, 8'd5, 8'd85, 8'd109, 8'd69, 8'd51, 8'd210, 8'd110, 8'd227, 8'd100, 8'd197, 8'd102, 8'd207, 8'd193, 8'd97, 8'd56, 8'd202, 8'd243, 8'd84, 8'd172, 8'd112, 8'd213, 8'd197, 8'd43, 8'd220, 8'd253, 8'd132, 8'd226, 8'd150, 8'd40, 8'd51, 8'd104, 8'd191, 8'd211, 8'd202, 8'd82, 8'd137, 8'd23, 8'd29, 8'd35, 8'd174, 8'd127, 8'd49, 8'd127, 8'd38, 8'd15, 8'd217, 8'd143, 8'd238, 8'd178, 8'd149, 8'd208, 8'd225, 8'd253, 8'd1, 8'd221, 8'd157, 8'd253, 8'd135, 8'd123, 8'd205, 8'd59, 8'd128, 8'd230, 8'd147, 8'd216, 8'd189, 8'd150, 8'd63, 8'd170, 8'd22, 8'd160, 8'd169, 8'd187, 8'd228, 8'd251, 8'd197, 8'd149, 8'd237, 8'd148, 8'd5, 8'd31, 8'd220, 8'd124, 8'd216, 8'd54, 8'd141, 8'd161, 8'd9, 8'd157, 8'd93, 8'd13, 8'd125, 8'd50, 8'd32, 8'd53, 8'd38, 8'd49, 8'd11, 8'd162, 8'd72, 8'd138, 8'd178, 8'd128, 8'd137, 8'd114, 8'd32, 8'd126, 8'd218, 8'd223, 8'd69, 8'd54, 8'd145, 8'd164, 8'd107, 8'd53, 8'd242, 8'd21, 8'd27, 8'd37, 8'd43, 8'd159, 8'd147, 8'd14, 8'd238, 8'd186, 8'd189, 8'd17, 8'd220, 8'd239, 8'd252, 8'd220, 8'd201, 8'd131, 8'd46, 8'd102, 8'd35, 8'd8, 8'd240, 8'd77, 8'd76, 8'd85, 8'd120, 8'd166, 8'd7, 8'd215, 8'd143, 8'd218, 8'd89, 8'd114, 8'd14, 8'd46, 8'd170, 8'd85, 8'd230, 8'd31, 8'd253, 8'd138, 8'd181, 8'd255, 8'd74, 8'd106, 8'd119, 8'd195, 8'd209, 8'd26, 8'd46, 8'd92, 8'd15, 8'd134, 8'd86, 8'd45, 8'd54, 8'd231, 8'd173, 8'd120, 8'd233, 8'd27, 8'd191, 8'd188, 8'd144, 8'd47, 8'd153, 8'd77, 8'd35, 8'd55, 8'd229, 8'd19, 8'd62, 8'd14, 8'd113, 8'd4, 8'd229, 8'd51, 8'd24, 8'd79, 8'd117, 8'd26, 8'd254, 8'd85, 8'd76, 8'd16, 8'd77, 8'd12, 8'd129, 8'd195, 8'd161, 8'd23, 8'd21, 8'd199, 8'd231, 8'd137, 8'd28, 8'd211 } ;
	// assign high value for square wave
	assign sqr_high = { 12'd2457, 12'd2866, 12'd3276, 12'd3686, 12'd4095 } ;
	// assign low value for square wave
	assign sqr_low = { 12'd1638, 12'd1228, 12'd819, 12'd410, 12'd0 } ; 

	// configure s2 as on/off switch
	always_ff @( negedge s2 )
		if ( ~s2 )
			onOff <= ~onOff ;

	always_comb begin
		// update data only when onOff enabled, otherwise default to 0V output data
		if ( onOff ) begin 
			if ( shape == 3'd1 ) // square wave mode
				if ( index < 8'd127 )
					next_data = sqr_high[depth] ;
				else
					next_data = sqr_low[depth] ;
			else if ( shape == 3'd5 ) // sample & hold mode
				next_data = SnH_value ;
			else
				next_data = dataTable[index] ; // all other modes
		end else
			next_data = 12'd0 ; // off
	end

	always_ff @( posedge wclk, negedge reset_n ) begin
		if ( ~reset_n )
			{ data, index, SnH_value, SnH_index_2 } <= '0 ; // reset conditions
		else begin 
			data <= next_data ;
			index <= index + 1'b1 ;
			if ( { shape, index } == { 3'd5, 8'd0 } || { shape, index } == { 3'd5, 8'd127 } ) begin // sample & hold mode
				SnH_value <= dataTable[SnH_index[SnH_index_2]] ; // "randomly" select sample & hold value
				SnH_index_2 <= SnH_index_2 + 1'b1 ;
			end else
				SnH_value <= SnH_value ;
		end  
	end

endmodule
